-- ALU.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU_INTF IS
	PORT (
		OPCODE_BUS : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		MUX_OUT_BUS : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ACC_DATA_OUT_BUS : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		OUTPUT_BUS : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ALU_INTF;

ARCHITECTURE ALU_ARCH OF ALU_INTF IS

BEGIN
	MAIN : PROCESS (OPCODE_BUS, MUX_OUT_BUS, ACC_DATA_OUT_BUS)
		VARIABLE A : unsigned(7 DOWNTO 0);
		VARIABLE B : unsigned(7 DOWNTO 0);
		VARIABLE TMP16 : unsigned (15 DOWNTO 0);
	BEGIN
		A := unsigned(ACC_DATA_OUT_BUS);
		B := unsigned(MUX_OUT_BUS);

		CASE(OPCODE_BUS) IS
			WHEN "000" =>
			OUTPUT_BUS <= STD_LOGIC_VECTOR(A);
			WHEN "001" =>
			OUTPUT_BUS <= STD_LOGIC_VECTOR(b);
			WHEN "010" =>
			TMP16 := A * B;
			OUTPUT_BUS <= STD_LOGIC_VECTOR(TMP16(7 DOWNTO 0));
			WHEN "011" =>
			OUTPUT_BUS <= STD_LOGIC_VECTOR(A SRL 1);
			WHEN "100" =>
			OUTPUT_BUS <= STD_LOGIC_VECTOR(A + B);
			WHEN OTHERS => OUTPUT_BUS <= "00000000";
		END CASE;
	END PROCESS MAIN;

END ALU_ARCH;