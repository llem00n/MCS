-- MUX.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_INTF IS
	PORT (
		SELECT_IN : IN STD_LOGIC;
		RAM_DATA_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		DATA_IN_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END MUX_INTF;

ARCHITECTURE MUX_ARCH OF MUX_INTF IS
	SIGNAL DEFAULT_VAL : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	DEFAULT_VAL <= "00000000";

	MAIN : PROCESS (SELECT_IN, DATA_IN_BUS, RAM_DATA_BUS)
	BEGIN
		CASE (SELECT_IN) IS
			WHEN '0' =>
				DATA_OUT <= DATA_IN_BUS;
			WHEN '1' =>
				DATA_OUT <= RAM_DATA_BUS;
			WHEN OTHERS =>
				DATA_OUT <= DEFAULT_VAL;
		END CASE;
	END PROCESS MAIN;
END MUX_ARCH;