-- DECODER.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DECODER_INTF IS
	PORT (
		CLOCK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		ACC_DATA_OUT_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		COMM_ONES : OUT STD_LOGIC;
		COMM_DECS : OUT STD_LOGIC;
		COMM_HUNDREDS : OUT STD_LOGIC;
		SEG_A : OUT STD_LOGIC;
		SEG_B : OUT STD_LOGIC;
		SEG_C : OUT STD_LOGIC;
		SEG_D : OUT STD_LOGIC;
		SEG_E : OUT STD_LOGIC;
		SEG_F : OUT STD_LOGIC;
		SEG_G : OUT STD_LOGIC;
		DP : OUT STD_LOGIC);
END DECODER_INTF;

ARCHITECTURE DECODER_ARCH OF DECODER_INTF IS
	SIGNAL ONES_BUS : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	SIGNAL DECS_BUS : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
	SIGNAL HONDREDS_BUS : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";

BEGIN
	BIN_TO_BCD : PROCESS (ACC_DATA_OUT_BUS)
		VARIABLE hex_src : STD_LOGIC_VECTOR(7 DOWNTO 0);
		VARIABLE bcd : STD_LOGIC_VECTOR(11 DOWNTO 0);
	BEGIN
		bcd := (OTHERS => '0');
		hex_src := ACC_DATA_OUT_BUS;

		FOR X IN hex_src'RANGE LOOP
			IF bcd(3 DOWNTO 0) > "0100" THEN
				bcd(3 DOWNTO 0) := bcd(3 DOWNTO 0) + "0011";
			END IF;
			IF bcd(7 DOWNTO 4) > "0100" THEN
				bcd(7 DOWNTO 4) := bcd(7 DOWNTO 4) + "0011";
			END IF;
			IF bcd(11 DOWNTO 8) > "0100" THEN
				bcd(11 DOWNTO 8) := bcd(11 DOWNTO 8) + "0011";
			END IF;

			bcd := bcd(10 DOWNTO 0) & hex_src(hex_src'left);
			hex_src := hex_src(hex_src'left - 1 DOWNTO hex_src'right) & '0';
		END LOOP;

		HONDREDS_BUS <= bcd (11 DOWNTO 8);
		DECS_BUS <= bcd (7 DOWNTO 4);
		ONES_BUS <= bcd (3 DOWNTO 0);

	END PROCESS BIN_TO_BCD;

	INDICATE : PROCESS (CLOCK)
		TYPE DIGIT_TYPE IS (ONES, DECS, HUNDREDS);

		VARIABLE CUR_DIGIT : DIGIT_TYPE := ONES;
		VARIABLE DIGIT_VAL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
		VARIABLE DIGIT_CTRL : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
		VARIABLE COMMONS_CTRL : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";

	BEGIN
		IF (rising_edge(CLOCK)) THEN
			IF (RESET = '0') THEN
				CASE CUR_DIGIT IS
					WHEN ONES =>
						DIGIT_VAL := ONES_BUS;
						CUR_DIGIT := DECS;
						COMMONS_CTRL := "001";
					WHEN DECS =>
						DIGIT_VAL := DECS_BUS;
						CUR_DIGIT := HUNDREDS;
						COMMONS_CTRL := "010";
					WHEN HUNDREDS =>
						DIGIT_VAL := HONDREDS_BUS;
						CUR_DIGIT := ONES;
						COMMONS_CTRL := "100";
					WHEN OTHERS =>
						DIGIT_VAL := ONES_BUS;
						CUR_DIGIT := ONES;
						COMMONS_CTRL := "000";
				END CASE;

				CASE DIGIT_VAL IS
					WHEN "0000" => DIGIT_CTRL := "1111110";
					WHEN "0001" => DIGIT_CTRL := "0110000";
					WHEN "0010" => DIGIT_CTRL := "1101101";
					WHEN "0011" => DIGIT_CTRL := "1111001";
					WHEN "0100" => DIGIT_CTRL := "0110011";
					WHEN "0101" => DIGIT_CTRL := "1011011";
					WHEN "0110" => DIGIT_CTRL := "1011111";
					WHEN "0111" => DIGIT_CTRL := "1110000";
					WHEN "1000" => DIGIT_CTRL := "1111111";
					WHEN "1001" => DIGIT_CTRL := "1111011";
					WHEN OTHERS => DIGIT_CTRL := "0000000";
				END CASE;
			ELSE
				DIGIT_VAL := ONES_BUS;
				CUR_DIGIT := ONES;
				COMMONS_CTRL := "000";
			END IF;

			COMM_ONES <= COMMONS_CTRL(0);
			COMM_DECS <= COMMONS_CTRL(1);
			COMM_HUNDREDS <= COMMONS_CTRL(2);

			SEG_A <= DIGIT_CTRL(6);
			SEG_B <= DIGIT_CTRL(5);
			SEG_C <= DIGIT_CTRL(4);
			SEG_D <= DIGIT_CTRL(3);
			SEG_E <= DIGIT_CTRL(2);
			SEG_F <= DIGIT_CTRL(1);
			SEG_G <= DIGIT_CTRL(0);
			DP <= '0';

		END IF;
	END PROCESS INDICATE;

END DECODER_ARCH;