-- ALU.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU_INTF IS
	PORT (
		OP_CODE_BUS : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		MUX_OUT_BUS : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ACC_DATA_OUT_BUS : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ACC_DATA_IN_BUS : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ALU_INTF;

ARCHITECTURE ALU_ARCH OF ALU_INTF IS

BEGIN
	ALU : PROCESS (OP_CODE_BUS, MUX_OUT_BUS, ACC_DATA_OUT_BUS)
		VARIABLE A : unsigned(7 DOWNTO 0);
		VARIABLE B : unsigned(7 DOWNTO 0);
		VARIABLE TEMP_MUL : unsigned (15 DOWNTO 0);
	BEGIN
		A := unsigned(ACC_DATA_OUT_BUS);
		B := unsigned(MUX_OUT_BUS);

		CASE(OP_CODE_BUS) IS
			WHEN "00" => ACC_DATA_IN_BUS <= STD_LOGIC_VECTOR(B);
			WHEN "01" => TEMP_MUL := (A * B);
			ACC_DATA_IN_BUS <= STD_LOGIC_VECTOR(TEMP_MUL(7 DOWNTO 0));
			WHEN "10" => ACC_DATA_IN_BUS <= STD_LOGIC_VECTOR(A SRL 1);
			WHEN "11" => ACC_DATA_IN_BUS <= STD_LOGIC_VECTOR(A + B);
			WHEN OTHERS => ACC_DATA_IN_BUS <= "00000000";
		END CASE;
	END PROCESS ALU;

END ALU_ARCH;