-- ACC.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ACC_INTF IS
	PORT (
		CLOCK : IN STD_LOGIC;
		DATA_IN_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		WR : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		DATA_OUT_BUS : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END ACC_INTF;

ARCHITECTURE ACC_ARCH OF ACC_INTF IS
	SIGNAL DATA : STD_LOGIC_VECTOR (7 DOWNTO 0);
BEGIN
	MAIN : PROCESS (CLOCK, DATA)
	BEGIN
		IF (rising_edge(CLOCK)) THEN
			IF (RST = '1') THEN
				DATA <= "00000000";
			ELSIF (WR = '1') THEN
				DATA <= DATA_IN_BUS;
			END IF;
		END IF;
		
		DATA_OUT_BUS <= DATA;
	END PROCESS MAIN;

END ACC_ARCH;