-- RAM.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RAM_INTF IS
	PORT (
		CLOCK : IN STD_LOGIC;
		WR : IN STD_LOGIC;
		DATA_IN_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		ADDRESS_BUS : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END RAM_INTF;

ARCHITECTURE RAM_ARCH OF RAM_INTF IS
	TYPE ram_type IS ARRAY (3 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RAM_UNIT : ram_type := (OTHERS => (OTHERS => '0'));
BEGIN
	RAM_IN : PROCESS (CLOCK)
	BEGIN
		IF (rising_edge(CLOCK)) THEN
			IF (WR = '1') THEN
				RAM_UNIT(conv_integer(ADDRESS_BUS)) <= DATA_IN_BUS;
			END IF;
		END IF;
	END PROCESS RAM_IN;
	
	RAM_OUT : PROCESS (CLOCK)
	BEGIN
		IF (rising_edge(CLOCK)) THEN
			DATA_OUT <= RAM_UNIT(conv_integer(ADDRESS_BUS));
		END IF;
	END PROCESS RAM_OUT;
END RAM_ARCH;