-- MUX.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_INTF IS
	PORT (
		SEL_IN_BUS : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		RAM_DATA_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		DATA_INPUT_BUS : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END MUX_INTF;

ARCHITECTURE MUX_ARCH OF MUX_INTF IS
	SIGNAL CONST : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	CONST <= "00000000";
	MUX : PROCESS (SEL_IN_BUS, DATA_INPUT_BUS, RAM_DATA_BUS)
	BEGIN
		CASE (SEL_IN_BUS) IS
			WHEN "00" => DATA_OUT <= DATA_INPUT_BUS;
			WHEN "01" => DATA_OUT <= RAM_DATA_BUS;
			WHEN OTHERS => DATA_OUT <= CONST;
		END CASE;
	END PROCESS;
END MUX_ARCH;